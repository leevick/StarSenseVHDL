library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top is

end top;

architecture Behavioral of top is

begin


end Behavioral;

